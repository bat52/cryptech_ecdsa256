/* Values from "Suite B Implementer's Guide to FIPS 186-3 (ECDSA)" */

localparam [255:0] ECDSA_P256_D_NSA =
	{32'h70a12c2d, 32'hb16845ed, 32'h56ff68cf, 32'hc21a472b,
	 32'h3f04d7d6, 32'h851bf634, 32'h9f2d7d5b, 32'h3452b38a};

localparam [255:0] ECDSA_P256_QX_NSA =
	{32'h8101ece4, 32'h7464a6ea, 32'hd70cf69a, 32'h6e2bd3d8,
	 32'h8691a326, 32'h2d22cba4, 32'hf7635eaf, 32'hf26680a8};
	 
localparam [255:0] ECDSA_P256_QY_NSA =
	{32'hd8a12ba6, 32'h1d599235, 32'hf67d9cb4, 32'hd58f1783,
	 32'hd3ca43e7, 32'h8f0a5aba, 32'ha6240799, 32'h36c0c3a9};
	 
localparam [255:0] ECDSA_P256_K_NSA =
	{32'h580ec00d, 32'h85643433, 32'h4cef3f71, 32'hecaed496,
	 32'h5b12ae37, 32'hfa47055b, 32'h1965c7b1, 32'h34ee45d0};

localparam [255:0] ECDSA_P256_RX_NSA =
	{32'h7214bc96, 32'h47160bbd, 32'h39ff2f80, 32'h533f5dc6,
	 32'hddd70ddf, 32'h86bb8156, 32'h61e805d5, 32'hd4e6f27c};
	 
localparam [255:0] ECDSA_P256_RY_NSA =
	{32'h8b81e3e9, 32'h77597110, 32'hc7cf2633, 32'h435b2294,
	 32'hb7264298, 32'h7defd3d4, 32'h007e1cfc, 32'h5df84541};

